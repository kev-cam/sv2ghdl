// Simple 2-input OR gate
module or_gate (
    input a,
    input b,
    output y
);

or or1 (y, a, b);

endmodule
