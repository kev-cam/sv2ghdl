// Simple NOT gate (inverter)
module not_gate (
    input a,
    output y
);

not not1 (y, a);

endmodule
