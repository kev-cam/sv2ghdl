// Simple 2-input AND gate
module and_gate (
    input a,
    input b,
    output y
);

and and1 (y, a, b);

endmodule
