// Simple 2-input XOR gate
module xor_gate (
    input a,
    input b,
    output y
);

assign y = a ^ b;

endmodule
